module and_gate
(
    input w_a,
    input w_b,
    output y
);

assign y = w_a & w_b;

endmodule